module OR7 (
    input  a, b, c, d, e, f, g,
    output y
);
    assign y = a | b | c | d | e | f | g;
endmodule
