module OR9 (
    input  a, b, c, d, e, f, g, h, i,
    output y
);
    assign y = a | b | c | d | e | f | g | h | i;
endmodule
