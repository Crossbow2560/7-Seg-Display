module OR8 (
    input  a, b, c, d, e, f, g, h,
    output y
);
    assign y = a | b | c | d | e | f | g | h;
endmodule
